module tb();
  reg [3:0] a,b;
  reg cin;
  wire [3:0] s;
  wire c;
  //instanciate the design under test 
  fa
